`timescale 1ns / 1ps
`default_nettype none

module top_level();
  graphics gr();
endmodule

`default_nettype wire